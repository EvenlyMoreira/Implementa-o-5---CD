LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY Cod6x3 IS
  PORT(
    A, B, C, D, E, F: IN STD_LOGIC;
    s: OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END ENTITY Cod6x3;

ARCHITECTURE log OF Cod6x3 IS
BEGIN
s(2) <=((NOT A) AND (NOT B) AND (NOT C) AND (NOT D));
s(1) <=((NOT A) AND (NOT B) AND (NOT E) AND (NOT F)) OR ((NOT A) AND (NOT B) AND D) OR ((NOT A) AND (NOT B) AND C);
s(0) <=((NOT A) AND (NOT C) AND (NOT E) AND F) OR ((NOT A) AND (NOT C) AND D) OR ((NOT A) AND B);
END ARCHITECTURE log;
